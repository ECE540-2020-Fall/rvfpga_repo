FFFE0E1300010E37
408E8E9380001EB7
800015B701CEA023
0005A28340058593
4045051380001537
005520230102D293
00000000FE0002E3
